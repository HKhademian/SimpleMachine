module Computer(
	ResetN, Clock, ABCD
    );


endmodule
